-- lab3.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lab3 is
	port (
		clk_clk                               : in    std_logic                    := '0'; --                            clk.clk
		opencores_i2c_0_export_0_scl_pad_io   : inout std_logic                    := '0'; --       opencores_i2c_0_export_0.scl_pad_io
		opencores_i2c_0_export_0_sda_pad_io   : inout std_logic                    := '0'; --                               .sda_pad_io
		pio_0_external_connection_export      : out   std_logic_vector(3 downto 0);        --      pio_0_external_connection.export
		pio_1_external_connection_export      : out   std_logic_vector(3 downto 0);        --      pio_1_external_connection.export
		pio_2_external_connection_export      : out   std_logic_vector(3 downto 0);        --      pio_2_external_connection.export
		pio_3_external_connection_export      : out   std_logic_vector(3 downto 0);        --      pio_3_external_connection.export
		pio_bouton_external_connection_export : in    std_logic                    := '0'; -- pio_bouton_external_connection.export
		reset_reset_n                         : in    std_logic                    := '0'  --                          reset.reset_n
	);
end entity lab3;

architecture rtl of lab3 is	
	component lab3 is
		port (
			clk_clk                               : in    std_logic                    := 'X'; -- clk
			opencores_i2c_0_export_0_scl_pad_io   : inout std_logic                    := 'X'; -- scl_pad_io
			opencores_i2c_0_export_0_sda_pad_io   : inout std_logic                    := 'X'; -- sda_pad_io
			pio_0_external_connection_export      : out   std_logic_vector(3 downto 0);        -- export
			pio_1_external_connection_export      : out   std_logic_vector(3 downto 0);        -- export
			pio_2_external_connection_export      : out   std_logic_vector(3 downto 0);        -- export
			pio_3_external_connection_export      : out   std_logic_vector(3 downto 0);        -- export
			reset_reset_n                         : in    std_logic                    := 'X'; -- reset_n
			pio_bouton_external_connection_export : in    std_logic                    := 'X'  -- export
		);
	end component lab3;
begin
	u0 : component lab3
		port map (
			clk_clk                               => CONNECTED_TO_clk_clk,                               --                            clk.clk
			opencores_i2c_0_export_0_scl_pad_io   => CONNECTED_TO_opencores_i2c_0_export_0_scl_pad_io,   --       opencores_i2c_0_export_0.scl_pad_io
			opencores_i2c_0_export_0_sda_pad_io   => CONNECTED_TO_opencores_i2c_0_export_0_sda_pad_io,   --                               .sda_pad_io
			pio_0_external_connection_export      => CONNECTED_TO_pio_0_external_connection_export,      --      pio_0_external_connection.export
			pio_1_external_connection_export      => CONNECTED_TO_pio_1_external_connection_export,      --      pio_1_external_connection.export
			pio_2_external_connection_export      => CONNECTED_TO_pio_2_external_connection_export,      --      pio_2_external_connection.export
			pio_3_external_connection_export      => CONNECTED_TO_pio_3_external_connection_export,      --      pio_3_external_connection.export
			reset_reset_n                         => CONNECTED_TO_reset_reset_n,                         --                          reset.reset_n
			pio_bouton_external_connection_export => CONNECTED_TO_pio_bouton_external_connection_export  -- pio_bouton_external_connection.export
		);

